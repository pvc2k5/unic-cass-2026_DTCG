* NGSPICE file created from user_project_wrapper.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_Filler400 abstract view
.subckt sg13g2_Filler400 iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_IOPadOut30mA abstract view
.subckt sg13g2_IOPadOut30mA c2p iovdd iovss pad vdd vss
.ends

* Black-box entry subcircuit for bondpad_70x70 abstract view
.subckt bondpad_70x70 pad
.ends

* Black-box entry subcircuit for sg13g2_Filler4000 abstract view
.subckt sg13g2_Filler4000 iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_IOPadIOVdd abstract view
.subckt sg13g2_IOPadIOVdd iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_IOPadIn abstract view
.subckt sg13g2_IOPadIn iovdd iovss p2c pad vdd vss
.ends

* Black-box entry subcircuit for sg13g2_Filler1000 abstract view
.subckt sg13g2_Filler1000 iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_IOPadVdd abstract view
.subckt sg13g2_IOPadVdd iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_IOPadIOVss abstract view
.subckt sg13g2_IOPadIOVss iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_IOPadVss abstract view
.subckt sg13g2_IOPadVss iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_Corner abstract view
.subckt sg13g2_Corner iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_Filler200 abstract view
.subckt sg13g2_Filler200 iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_IOPadAnalog abstract view
.subckt sg13g2_IOPadAnalog iovdd iovss pad padres vdd vss
.ends

.subckt user_project_wrapper IOVDD IOVSS VDD VSS analog_io_0 analog_io_1 io_clock_PAD
+ io_reset_PAD ui_PAD[0] ui_PAD[10] ui_PAD[11] ui_PAD[12] ui_PAD[13] ui_PAD[14] ui_PAD[15]
+ ui_PAD[1] ui_PAD[2] ui_PAD[3] ui_PAD[4] ui_PAD[5] ui_PAD[6] ui_PAD[7] ui_PAD[8]
+ ui_PAD[9] uo_PAD[0] uo_PAD[10] uo_PAD[11] uo_PAD[12] uo_PAD[13] uo_PAD[14] uo_PAD[15]
+ uo_PAD[1] uo_PAD[2] uo_PAD[3] uo_PAD[4] uo_PAD[5] uo_PAD[6] uo_PAD[7] uo_PAD[8]
+ uo_PAD[9]
XIO_FILL_IO_NORTH_1_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
Xsg13g2_IOPadOut30mA_uo\[9\].uo sg13g2_IOPadOut30mA_uo\[9\].uo/c2p IOVDD IOVSS uo_PAD[9]
+ VDD VSS sg13g2_IOPadOut30mA
XIO_FILL_IO_NORTH_4_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_BOND_sg13g2_IOPadIn_ui\[7\].ui ui_PAD[7] bondpad_70x70
XIO_FILL_IO_SOUTH_3_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
Xsg13g2_IOPadIOVdd_south IOVDD IOVSS VDD VSS sg13g2_IOPadIOVdd
XIO_FILL_IO_NORTH_7_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_NORTH_0_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_BOND_sg13g2_IOPadIn_ui\[14\].ui ui_PAD[14] bondpad_70x70
XIO_FILL_IO_EAST_12_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_SOUTH_1_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_BOND_sg13g2_IOPadOut30mA_uo\[14\].uo uo_PAD[14] bondpad_70x70
Xsg13g2_IOPadIn_ui\[7\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[7\].ui/p2c ui_PAD[7] VDD
+ VSS sg13g2_IOPadIn
XIO_FILL_IO_SOUTH_4_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_WEST_11_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
Xsg13g2_IOPad_io_clock IOVDD IOVSS sg13g2_IOPad_io_clock/p2c io_clock_PAD VDD VSS
+ sg13g2_IOPadIn
XIO_FILL_IO_WEST_2_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_SOUTH_7_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_NORTH_10_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
Xsg13g2_IOPadIn_ui\[11\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[11\].ui/p2c ui_PAD[11]
+ VDD VSS sg13g2_IOPadIn
XIO_FILL_IO_EAST_0_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_BOND_sg13g2_IOPadVss_west VSS bondpad_70x70
XIO_FILL_IO_NORTH_13_20 IOVDD IOVSS VDD VSS sg13g2_Filler1000
Xsg13g2_IOPad_io_reset IOVDD IOVSS sg13g2_IOPad_io_reset/p2c io_reset_PAD VDD VSS
+ sg13g2_IOPadIn
XIO_FILL_IO_SOUTH_1_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_SOUTH_10_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_SOUTH_13_20 IOVDD IOVSS VDD VSS sg13g2_Filler1000
XIO_FILL_IO_EAST_10_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_EAST_10_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_NORTH_9_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_EAST_2_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_EAST_13_20 IOVDD IOVSS VDD VSS sg13g2_Filler1000
XIO_FILL_IO_WEST_12_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_BOND_sg13g2_IOPadOut30mA_uo\[2\].uo uo_PAD[2] bondpad_70x70
Xsg13g2_IOPadVdd_south IOVDD IOVSS VDD VSS sg13g2_IOPadVdd
XIO_FILL_IO_EAST_5_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_WEST_0_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
Xsg13g2_IOPadOut30mA_uo\[2\].uo sg13g2_IOPadOut30mA_uo\[2\].uo/c2p IOVDD IOVSS uo_PAD[2]
+ VDD VSS sg13g2_IOPadOut30mA
Xsg13g2_IOPadIn_ui\[14\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[14\].ui/p2c ui_PAD[14]
+ VDD VSS sg13g2_IOPadIn
Xsg13g2_IOPadIOVss_south IOVDD IOVSS VDD VSS sg13g2_IOPadIOVss
XIO_BOND_sg13g2_IOPadVss_east VSS bondpad_70x70
XIO_FILL_IO_EAST_8_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_BOND_sg13g2_IOPadIn_ui\[0\].ui ui_PAD[0] bondpad_70x70
Xsg13g2_IOPadVss_west IOVDD IOVSS VDD VSS sg13g2_IOPadVss
XIO_CORNER_NORTH_EAST_INST IOVDD IOVSS VDD VSS sg13g2_Corner
XIO_FILL_IO_EAST_9_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
Xsg13g2_IOPadIOVdd_north IOVDD IOVSS VDD VSS sg13g2_IOPadIOVdd
Xsg13g2_IOPadOut30mA_uo\[11\].uo sg13g2_IOPadOut30mA_uo\[11\].uo/c2p IOVDD IOVSS uo_PAD[11]
+ VDD VSS sg13g2_IOPadOut30mA
Xsg13g2_IOPadIn_ui\[0\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[0\].ui/p2c ui_PAD[0] VDD
+ VSS sg13g2_IOPadIn
XIO_FILL_IO_NORTH_7_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_BOND_sg13g2_IOPadOut30mA_uo\[5\].uo uo_PAD[5] bondpad_70x70
XIO_FILL_IO_WEST_10_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_NORTH_12_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_NORTH_13_25 IOVDD IOVSS VDD VSS sg13g2_Filler400
Xsg13g2_IOPadOut30mA_uo\[5\].uo sg13g2_IOPadOut30mA_uo\[5\].uo/c2p IOVDD IOVSS uo_PAD[5]
+ VDD VSS sg13g2_IOPadOut30mA
XIO_FILL_IO_WEST_2_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
Xsg13g2_IOPadVss_east IOVDD IOVSS VDD VSS sg13g2_IOPadVss
XIO_BOND_sg13g2_IOPadIn_ui\[3\].ui ui_PAD[3] bondpad_70x70
XIO_FILL_IO_WEST_9_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_WEST_5_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_SOUTH_13_25 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_BOND_sg13g2_IOPadVdd_west VDD bondpad_70x70
Xsg13g2_IOPadOut30mA_uo\[14\].uo sg13g2_IOPadOut30mA_uo\[14\].uo/c2p IOVDD IOVSS uo_PAD[14]
+ VDD VSS sg13g2_IOPadOut30mA
XIO_BOND_sg13g2_IOPadIn_ui\[10\].ui ui_PAD[10] bondpad_70x70
XIO_FILL_IO_EAST_7_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_CORNER_SOUTH_EAST_INST IOVDD IOVSS VDD VSS sg13g2_Corner
XIO_BOND_sg13g2_IOPadOut30mA_uo\[10\].uo uo_PAD[10] bondpad_70x70
XIO_FILL_IO_WEST_8_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
Xsg13g2_IOPadIn_ui\[3\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[3\].ui/p2c ui_PAD[3] VDD
+ VSS sg13g2_IOPadIn
XIO_FILL_IO_SOUTH_12_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_EAST_13_25 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_NORTH_13_27 IOVDD IOVSS VDD VSS sg13g2_Filler200
XIO_CORNER_NORTH_WEST_INST IOVDD IOVSS VDD VSS sg13g2_Corner
XIO_BOND_sg13g2_IOPadOut30mA_uo\[8\].uo uo_PAD[8] bondpad_70x70
Xsg13g2_IOPadVss_south IOVDD IOVSS VDD VSS sg13g2_IOPadVss
XIO_FILL_IO_SOUTH_8_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_NORTH_5_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_SOUTH_13_27 IOVDD IOVSS VDD VSS sg13g2_Filler200
Xsg13g2_IOPadVdd_north IOVDD IOVSS VDD VSS sg13g2_IOPadIOVdd
Xsg13g2_IOPadOut30mA_uo\[8\].uo sg13g2_IOPadOut30mA_uo\[8\].uo/c2p IOVDD IOVSS uo_PAD[8]
+ VDD VSS sg13g2_IOPadOut30mA
XIO_FILL_IO_NORTH_10_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_BOND_sg13g2_IOPadIn_ui\[6\].ui ui_PAD[6] bondpad_70x70
XIO_BOND_sg13g2_IOPadVdd_east VDD bondpad_70x70
Xsg13g2_IOPadIOVss_north IOVDD IOVSS VDD VSS sg13g2_IOPadIOVss
XIO_FILL_IO_NORTH_2_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_BOND_sg13g2_IOPadIn_ui\[13\].ui ui_PAD[13] bondpad_70x70
Xsg13g2_IOPadVdd_west IOVDD IOVSS VDD VSS sg13g2_IOPadVdd
XIO_FILL_IO_EAST_13_27 IOVDD IOVSS VDD VSS sg13g2_Filler200
XIO_FILL_IO_WEST_7_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_BOND_sg13g2_IOPadOut30mA_uo\[13\].uo uo_PAD[13] bondpad_70x70
XIO_FILL_IO_NORTH_5_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
Xsg13g2_IOPadIn_ui\[6\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[6\].ui/p2c ui_PAD[6] VDD
+ VSS sg13g2_IOPadIn
XIO_FILL_IO_EAST_5_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_SOUTH_10_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_NORTH_8_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_SOUTH_2_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_CORNER_SOUTH_WEST_INST IOVDD IOVSS VDD VSS sg13g2_Corner
XIO_FILL_IO_SOUTH_6_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_SOUTH_5_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_NORTH_3_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_WEST_12_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_BOND_sg13g2_IOPadIn_ui\[9\].ui ui_PAD[9] bondpad_70x70
Xsg13g2_IOPadIn_ui\[10\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[10\].ui/p2c ui_PAD[10]
+ VDD VSS sg13g2_IOPadIn
Xsg13g2_IOPad_analog_io_0 IOVDD IOVSS analog_io_0 sg13g2_IOPad_analog_io_0/padres
+ VDD VSS sg13g2_IOPadAnalog
Xsg13g2_IOPadVdd_east IOVDD IOVSS VDD VSS sg13g2_IOPadVdd
XIO_FILL_IO_SOUTH_8_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_NORTH_11_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
Xsg13g2_IOPad_analog_io_1 IOVDD IOVSS analog_io_1 sg13g2_IOPad_analog_io_1/padres
+ VDD VSS sg13g2_IOPadAnalog
XIO_FILL_IO_WEST_5_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
Xsg13g2_IOPadIn_ui\[9\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[9\].ui/p2c ui_PAD[9] VDD
+ VSS sg13g2_IOPadIn
XIO_FILL_IO_SOUTH_11_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_EAST_3_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_BOND_sg13g2_IOPad_analog_io_0 analog_io_0 bondpad_70x70
XIO_FILL_IO_EAST_0_20 IOVDD IOVSS VDD VSS sg13g2_Filler1000
Xsg13g2_IOPadVss_north IOVDD IOVSS VDD VSS sg13g2_IOPadIOVss
XIO_BOND_sg13g2_IOPadOut30mA_uo\[1\].uo uo_PAD[1] bondpad_70x70
XIO_FILL_IO_EAST_11_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_SOUTH_4_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
Xsg13g2_IOPadIn_ui\[13\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[13\].ui/p2c ui_PAD[13]
+ VDD VSS sg13g2_IOPadIn
XIO_BOND_sg13g2_IOPad_io_clock io_clock_PAD bondpad_70x70
Xsg13g2_IOPadOut30mA_uo\[1\].uo sg13g2_IOPadOut30mA_uo\[1\].uo/c2p IOVDD IOVSS uo_PAD[1]
+ VDD VSS sg13g2_IOPadOut30mA
XIO_FILL_IO_EAST_3_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_BOND_sg13g2_IOPad_analog_io_1 analog_io_1 bondpad_70x70
XIO_FILL_IO_EAST_13_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_NORTH_1_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_EAST_6_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
Xsg13g2_IOPadOut30mA_uo\[10\].uo sg13g2_IOPadOut30mA_uo\[10\].uo/c2p IOVDD IOVSS uo_PAD[10]
+ VDD VSS sg13g2_IOPadOut30mA
XIO_BOND_sg13g2_IOPad_io_reset io_reset_PAD bondpad_70x70
XIO_FILL_IO_EAST_9_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_BOND_sg13g2_IOPadIOVdd_south IOVDD bondpad_70x70
XIO_FILL_IO_WEST_3_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_BOND_sg13g2_IOPadOut30mA_uo\[4\].uo uo_PAD[4] bondpad_70x70
XIO_FILL_IO_EAST_1_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
Xsg13g2_IOPadOut30mA_uo\[4\].uo sg13g2_IOPadOut30mA_uo\[4\].uo/c2p IOVDD IOVSS uo_PAD[4]
+ VDD VSS sg13g2_IOPadOut30mA
XIO_BOND_sg13g2_IOPadVdd_south VDD bondpad_70x70
XIO_FILL_IO_SOUTH_2_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_WEST_0_20 IOVDD IOVSS VDD VSS sg13g2_Filler1000
XIO_BOND_sg13g2_IOPadIn_ui\[2\].ui ui_PAD[2] bondpad_70x70
Xsg13g2_IOPadOut30mA_uo\[13\].uo sg13g2_IOPadOut30mA_uo\[13\].uo/c2p IOVDD IOVSS uo_PAD[13]
+ VDD VSS sg13g2_IOPadOut30mA
XIO_FILL_IO_EAST_11_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_WEST_3_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
Xsg13g2_IOPadIn_ui\[2\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[2\].ui/p2c ui_PAD[2] VDD
+ VSS sg13g2_IOPadIn
XIO_FILL_IO_EAST_0_25 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_WEST_13_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_WEST_6_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_BOND_sg13g2_IOPadOut30mA_uo\[7\].uo uo_PAD[7] bondpad_70x70
XIO_FILL_IO_WEST_1_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_WEST_9_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
Xsg13g2_IOPadOut30mA_uo\[7\].uo sg13g2_IOPadOut30mA_uo\[7\].uo/c2p IOVDD IOVSS uo_PAD[7]
+ VDD VSS sg13g2_IOPadOut30mA
XIO_BOND_sg13g2_IOPadIn_ui\[5\].ui ui_PAD[5] bondpad_70x70
Xsg13g2_IOPadIOVss_west IOVDD IOVSS VDD VSS sg13g2_IOPadIOVss
XIO_FILL_IO_SOUTH_0_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_BOND_sg13g2_IOPadIn_ui\[12\].ui ui_PAD[12] bondpad_70x70
XIO_FILL_IO_EAST_0_27 IOVDD IOVSS VDD VSS sg13g2_Filler200
XIO_FILL_IO_NORTH_0_20 IOVDD IOVSS VDD VSS sg13g2_Filler1000
XIO_BOND_sg13g2_IOPadOut30mA_uo\[12\].uo uo_PAD[12] bondpad_70x70
Xsg13g2_IOPadIn_ui\[5\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[5\].ui/p2c ui_PAD[5] VDD
+ VSS sg13g2_IOPadIn
XIO_BOND_sg13g2_IOPadIOVss_south IOVSS bondpad_70x70
XIO_FILL_IO_NORTH_8_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_NORTH_3_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_BOND_sg13g2_IOPadIOVdd_north IOVDD bondpad_70x70
XIO_FILL_IO_WEST_11_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_NORTH_13_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_NORTH_6_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_SOUTH_0_20 IOVDD IOVSS VDD VSS sg13g2_Filler1000
Xsg13g2_IOPadIOVss_east IOVDD IOVSS VDD VSS sg13g2_IOPadIOVss
XIO_BOND_sg13g2_IOPadVss_south VSS bondpad_70x70
XIO_FILL_IO_WEST_0_25 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_NORTH_9_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_BOND_sg13g2_IOPadIn_ui\[8\].ui ui_PAD[8] bondpad_70x70
XIO_FILL_IO_WEST_10_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_SOUTH_3_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_BOND_sg13g2_IOPadIn_ui\[15\].ui ui_PAD[15] bondpad_70x70
XIO_BOND_sg13g2_IOPadIOVss_west IOVSS bondpad_70x70
XIO_BOND_sg13g2_IOPadOut30mA_uo\[15\].uo uo_PAD[15] bondpad_70x70
XIO_BOND_sg13g2_IOPadVdd_north IOVDD bondpad_70x70
XIO_FILL_IO_WEST_13_20 IOVDD IOVSS VDD VSS sg13g2_Filler1000
Xsg13g2_IOPadIn_ui\[8\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[8\].ui/p2c ui_PAD[8] VDD
+ VSS sg13g2_IOPadIn
XIO_FILL_IO_EAST_8_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_SOUTH_6_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_SOUTH_13_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_SOUTH_9_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_SOUTH_9_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_WEST_0_27 IOVDD IOVSS VDD VSS sg13g2_Filler200
XIO_FILL_IO_NORTH_12_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_NORTH_6_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_BOND_sg13g2_IOPadOut30mA_uo\[0\].uo uo_PAD[0] bondpad_70x70
XIO_FILL_IO_NORTH_11_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
Xsg13g2_IOPadIn_ui\[12\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[12\].ui/p2c ui_PAD[12]
+ VDD VSS sg13g2_IOPadIn
XIO_FILL_IO_SOUTH_12_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
Xsg13g2_IOPadOut30mA_uo\[0\].uo sg13g2_IOPadOut30mA_uo\[0\].uo/c2p IOVDD IOVSS uo_PAD[0]
+ VDD VSS sg13g2_IOPadOut30mA
XIO_BOND_sg13g2_IOPadIOVss_east IOVSS bondpad_70x70
XIO_FILL_IO_NORTH_0_25 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_WEST_8_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_EAST_1_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_EAST_12_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
Xsg13g2_IOPadIOVdd_west IOVDD IOVSS VDD VSS sg13g2_IOPadIOVdd
XIO_FILL_IO_EAST_4_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_EAST_6_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_SOUTH_11_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_BOND_sg13g2_IOPadIOVss_north IOVSS bondpad_70x70
XIO_FILL_IO_EAST_7_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_SOUTH_0_25 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_SOUTH_7_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_BOND_sg13g2_IOPadOut30mA_uo\[3\].uo uo_PAD[3] bondpad_70x70
XIO_FILL_IO_NORTH_0_27 IOVDD IOVSS VDD VSS sg13g2_Filler200
XIO_FILL_IO_NORTH_4_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
Xsg13g2_IOPadOut30mA_uo\[3\].uo sg13g2_IOPadOut30mA_uo\[3\].uo/c2p IOVDD IOVSS uo_PAD[3]
+ VDD VSS sg13g2_IOPadOut30mA
Xsg13g2_IOPadIn_ui\[15\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[15\].ui/p2c ui_PAD[15]
+ VDD VSS sg13g2_IOPadIn
Xsg13g2_IOPadIOVdd_east IOVDD IOVSS VDD VSS sg13g2_IOPadIOVdd
XIO_BOND_sg13g2_IOPadIn_ui\[1\].ui ui_PAD[1] bondpad_70x70
XIO_BOND_sg13g2_IOPadVss_north IOVSS bondpad_70x70
XIO_FILL_IO_WEST_13_25 IOVDD IOVSS VDD VSS sg13g2_Filler400
Xsg13g2_IOPadOut30mA_uo\[12\].uo sg13g2_IOPadOut30mA_uo\[12\].uo/c2p IOVDD IOVSS uo_PAD[12]
+ VDD VSS sg13g2_IOPadOut30mA
XIO_BOND_sg13g2_IOPadIOVdd_west IOVDD bondpad_70x70
XIO_FILL_IO_WEST_6_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_SOUTH_0_27 IOVDD IOVSS VDD VSS sg13g2_Filler200
Xsg13g2_IOPadIn_ui\[1\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[1\].ui/p2c ui_PAD[1] VDD
+ VSS sg13g2_IOPadIn
XIO_FILL_IO_EAST_4_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_WEST_1_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_BOND_sg13g2_IOPadOut30mA_uo\[6\].uo uo_PAD[6] bondpad_70x70
XIO_FILL_IO_WEST_4_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_WEST_13_27 IOVDD IOVSS VDD VSS sg13g2_Filler200
Xsg13g2_IOPadOut30mA_uo\[6\].uo sg13g2_IOPadOut30mA_uo\[6\].uo/c2p IOVDD IOVSS uo_PAD[6]
+ VDD VSS sg13g2_IOPadOut30mA
XIO_FILL_IO_SOUTH_5_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_FILL_IO_WEST_7_20 IOVDD IOVSS VDD VSS sg13g2_Filler400
XIO_FILL_IO_NORTH_2_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_BOND_sg13g2_IOPadIn_ui\[4\].ui ui_PAD[4] bondpad_70x70
XIO_BOND_sg13g2_IOPadIOVdd_east IOVDD bondpad_70x70
XIO_BOND_sg13g2_IOPadIn_ui\[11\].ui ui_PAD[11] bondpad_70x70
Xsg13g2_IOPadOut30mA_uo\[15\].uo sg13g2_IOPadOut30mA_uo\[15\].uo/c2p IOVDD IOVSS uo_PAD[15]
+ VDD VSS sg13g2_IOPadOut30mA
XIO_BOND_sg13g2_IOPadOut30mA_uo\[11\].uo uo_PAD[11] bondpad_70x70
Xsg13g2_IOPadIn_ui\[4\].ui IOVDD IOVSS sg13g2_IOPadIn_ui\[4\].ui/p2c ui_PAD[4] VDD
+ VSS sg13g2_IOPadIn
XIO_FILL_IO_WEST_4_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
XIO_BOND_sg13g2_IOPadOut30mA_uo\[9\].uo uo_PAD[9] bondpad_70x70
XIO_FILL_IO_EAST_2_0 IOVDD IOVSS VDD VSS sg13g2_Filler4000
.ends

